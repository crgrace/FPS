// File Name: regfile_assign.sv
// Engineer:  Carl Grace (crgrace@lbl.gov)
// Description:  Code used in regfile.sv for assignment
//          
///////////////////////////////////////////////////////////////////

config_bits[LVDS_TRIGGER] <= 8'h07;
config_bits[LVDS_CONFIG] <= 8'h07;
config_bits[CML_DRIVER] <= 8'h07;
config_bits[PREAMP] <= 8'h07;
config_bits[VOLTAGE_FOLLOWER] <= 8'h07;
config_bits[IMONITOR] <= 8'h00;
config_bits[SPARE0] <= 8'h00;
config_bits[SPARE1] <= 8'h00;
config_bits[SPARE2] <= 8'h00;


